/* Transmitter */
/* Controller Module */

/* Controller module for the transmitter
which has 4 state: IDLE, LOAD, TRANS, and HOLD,
which indicates, respectively, the transmitter is idle, 
the transmitter loads the data, the transmitter is 
transmitting  the data, the transmitter is preparing
for the next idle state. The controller output
relative signals to control the other module of the transmitter */

module TransmitterController
(
	input			clk,
	input			rst,
	input			ena,
	input			start,
	input			bit_done,
	input			baud_full,
	input			baud_txir,
	output reg	shift,		// shift the shift register
	output reg	load,			// load data to the shift register
	output reg	inc,			// increment the bit counter
	output reg	ena_baud,	// enable the baud generator
	output reg 	ena_bit,		// enable the bit counter
	output reg 	ena_inv,		// enable the inverter
	output reg  clear_baud,
	output reg	clear_bit,
	output reg	clear_shift,
	output reg	clear_inv,
	output reg	done
);

parameter IDLE		= 2'b00;	// idle state, where data is ready to be transmitted
parameter LOAD 	= 2'b01;	// load state, where data is loaded
parameter TRANS	= 2'b11;	// transmitting state, where data is transmitted

reg [1:0] pstate, nstate;

always @(posedge clk)
begin
	pstate <= nstate;
end

always @(pstate, rst, ena, start, bit_done, baud_full, baud_txir)
begin
	shift			= 1'b0;
	load			= 1'b0;
	inc			= 1'b0;
	ena_baud		= 1'b0;
	ena_bit 		= 1'b0;
	ena_inv		= 1'b0;
	clear_baud	= 1'b0;
	clear_bit	= 1'b0;
	clear_shift	= 1'b0;
	clear_inv	= 1'b0;
	done			= 1'b0;
	nstate 		= pstate;		// defaultly keep the present state in loop
	
	if(!rst) begin
		clear_baud	= 1'b1;
		clear_bit	= 1'b1;
		clear_shift	= 1'b1;
		clear_inv 	= 1'b1;
		nstate 		= IDLE;
	end
	else if(ena) begin
		case(pstate)
			IDLE: begin
			clear_baud	= 1'b1;
			clear_bit	= 1'b1;

			if(start)
				nstate = LOAD;					// start to transmit when pushbutton is pressed
			end
			
			LOAD: begin
				load		= 1'b1;				// load the data to the shift register
				nstate	= TRANS;				// move to the TRANS state
			end

			TRANS: begin
				ena_baud	= 1'b1;				// enable the baud generator
				ena_bit  = 1'b1;				// enable the bit counter
				
				if(bit_done) begin			// when 10 bits of data is counted, a frame of data is completed transmitting
					done		= 1'b1;
					nstate 	= IDLE;			// move to the IDLE state
				end
				
				if(baud_txir)
					ena_inv = 1'b1;
				
				if(baud_full) begin			// shift and increment every baud tick
					shift = 1'b1;
					inc 	= 1'b1;
				end	
			end
		
			default begin
				nstate = IDLE;					// IDLE state by default
			end
		endcase
	end
end
endmodule
