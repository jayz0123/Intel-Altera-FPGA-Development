library verilog;
use verilog.vl_types.all;
entity ClockBlk_vlg_vec_tst is
end ClockBlk_vlg_vec_tst;
