library verilog;
use verilog.vl_types.all;
entity ClockBlk_vlg_sample_tst is
    port(
        inclk0          : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end ClockBlk_vlg_sample_tst;
