library verilog;
use verilog.vl_types.all;
entity MIPS_System_vlg_vec_tst is
end MIPS_System_vlg_vec_tst;
